~~~~~~~~~~~~~~~~~>Y~5Z!@'0\>C<]6]'5\!+\!<C6A2G:\=>Y~~~~~~~~~~~~~~~~~>Y_:Q!R!JsZ6V6^9&@6:V6V}@'W_<T:Pbg2_?^9^96]'Z'JsK<AT6GsZ >YssC<A':]#F'Z=C&Gai:]s@'W_<T:PE6P'\!bsW<D=G<ch>Yssss\&G#F'i<F' G7l?\4Z0l%V0G<A{f7\$]'\szh>YssV=WsK<AT6Gh>Y>YR!P;Z'V0G&A6V;R%Z<A2_s\5+\!l4V':@^91V4Z=>Yss\&G#F'osZ=C&Gb+\!:]#F'h>YV=Wsq6[2E:\!R?^9^9~~~~~~~~~~~~~~~~~^9~s@6P<]70\>C<]6]'5\!7V0\7V!gKb^9~~~~~~~~~~~~~~~~~^9?Z1A2A*:V6Vh>YF VsZ6V6 G7l?\4Z0lbe}R?_h>Y>YV=G:G*7V0\7V!lgKbsZ >YssC<A':]#F'i:]s@'W_<T:PE6P'\!`7\$]'\sz^9ssss<F'C&Gs	s\&Gs@'W_<T:PE6P'\!bsW<D=G<cz^9ss6]77V0\7V!lgKbh>Y>YR!P;Z'V0G&A6V;R%Z<A2_s\57V0\7V!lgKbsZ >YQ6T:]^9ss#A<P6@ :]#F'^9ss1V4Z=>YssssP2@6:]#F':@^9ssssss$[6]sccqns\&G#F'osccccccccq^9ssssss$[6]sccqns\&G#F'oscccccccbq^9ssssss$[6]scbqns\&G#F'osccccccccq^9ssssss$[6]scbqns\&G#F'osccccccbcq^9ssssss$[6]sccqns\&G#F'osccccccccq^9ssssss$[6]sccqns\&G#F'oscccccbccq^9ssssss$[6]scbqns\&G#F'osccccccccq^9ssssss$[6]scbqns\&G#F'osccccbcccq^9ssssss$[6]sbcqns\&G#F'osccccccccq^9ssssss$[6]sbcqns\&G#F'oscccbccccq^9ssssss$[6]sbbqns\&G#F'osccccccccq^9ssssss$[6]sbbqns\&G#F'osccbcccccq^9ssssss$[6]sbcqns\&G#F'osccccccccq^9ssssss$[6]sbcqns\&G#F'oscbccccccq^9ssssss$[6]sbbqns\&G#F'osccccccccq^9ssssss$[6]sbbqns\&G#F'osbcccccccq^9ssssss$[6]s\'[6A ns\&G#F'osccccccccq^9ssss6]70R Vh>YssV=WsC!\0V @h>YV=Wsq6[2E:\!R?^9^9~~~~~~~~~~~~~~~~~^9~s^2Z=0\>C<]6]'>Y~~~~~~~~~~~~~~~~~>Y_:Q!R!JsZ6V6^9&@6:V6V}@'W_<T:Pbg2_?^9^96]'Z'Js^2Z=:@^9ss#\!G{Z=C&GZ=C&Gs	sZ= G7l?\4Z0l%V0G<A{ sW<D=G<ch>YssssK<AV*i:]s@'W_<T:PE6P'\!bsW<D=G<ch>Yssss\&G#F'\&G#F's	s\&Gs@'W_<T:PE6P'\!bsW<D=G<cz^9ss6]7>R:]h>Y>YR!P;Z'V0G&A6V;R%Z<A2_s\5>R:]sZ >Y>Yss@:T=R?7V0\7V!W6P<W6Aa	s@'W_<T:PE6P'\!bsW<D=G<ch>YssP<^#\=V=GsK<AT6GsZ >YssssC<A':]#F'Z=C&Gai:]s@'W_<T:PE6P'\!bsW<D=G<ch>Yssssss\&G#F'i<F' G7l?\4Z0l%V0G<A{f7\$]'\szh>YssssV=WsP<^#\=V=Gh>YssP<^#\=V=GsW6P<W6A+e:@^9ssss#\!G{Z=C&Gs	sZ= G7l?\4Z0l%V0G<A{ sW<D=G<ch>Yssssss\&G#F'i<F' G7l?\4Z0l%V0G<A{f7\$]'\szh>YssssV=WsP<^#\=V=Gh>YssssssQ6T:]^9sssssssss	sW6P<W6A+e#\!Gs^2C{Z=C&GW6P<W6Abh>Yssssssssbi7V0\7V!lgKbsC<A'>R#:]#F'la7V0\7V!z^9sssssssss	sK<AT6GsC<A'>R#7V0\7V!K<AV*<F'C&Gbh>Yssssssss`i+\!l4V'#\!Gs^2C{W6P<W6Aa+\!x6J\&G#F'z^9^9ssss6]7V;R%Z<A2_h