>9UZA@GP\^C\]V]GU\AK\A\CVARGZ\]>9>9_ZQARAJZVVV>9F@VZVVV@GWl_\TZPlR__>9>9V]GZGJK\AlTVGZ@>9C\AGZ]CFGZ]CFG	Z]@GWl_\TZPlEVPG\AW\D]G\>9\FGCFG	\FG@GWl_\TZPlEVPG\AW\D]G\>9V]WK\AlTVG>9>9RAP[ZGVPGFAVqV[REZ\AR_\UK\AlTVGZ@>9QVTZ]>9\FGCFGZ]CFGK\AZ]CFG>9V]WqV[REZ\AR_>9>9>9@VP\]WP\^C\]V]GU\AWVP\WVAK>9>9_ZQARAJZVVV>9F@VZVVV@GWl_\TZPlR__>9>9V]GZGJWVP\WVAlKZ@>9C\AGZ]CFG	Z]@GWl_\TZPlEVPG\A W\D]G\>9\FGCFG	\FG@GWl_\TZPlEVPG\AW\D]G\>9V]WWVP\WVAlK>9>9RAP[ZGVPGFAVqV[REZ\AR_\UWVP\WVAlKZ@>9QVTZ]>9CA\PV@@Z]CFG>9QVTZ]>9PR@VZ]CFGZ@>9D[V]\FGCFG>9D[V]\FGCFG>9D[V]\FGCFG>9D[V]\FGCFG>9D[V]\FGCFG>9D[V]\FGCFG>9D[V]\FGCFG>9D[V]\FGCFG>9D[V]\FGCFG>9D[V]\FGCFG>9D[V]\FGCFG>9D[V]\FGCFG>9D[V]\FGCFG>9D[V]\FGCFG>9D[V]\FGCFG>9D[V]\FGCFG>9D[V]\G[VA@\FGCFG>9V]WPR@V>9V]WCA\PV@@>9V]WqV[REZ\AR_>9>9>9^RZ]P\^C\]V]G>9>9_ZQARAJZVVV>9F@VZVVV@GWl_\TZPlR__>9>9V]GZGJ^RZ]Z@>9C\AGZ]CFGlZ]CFGl	Z]@GWl_\TZPlEVPG\A W\D]G\>9K\AxVJ	Z]@GWl_\TZPlEVPG\AW\D]G\>9\FGCFG\FGCFG	\FG@GWl_\TZPlEVPG\AW\D]G\>9V]W^RZ]>9>9RAP[ZGVPGFAVqV[REZ\AR_\U^RZ]Z@>9>9@ZT]R_WVP\WVAWVP\WVA	@GWl_\TZPlEVPG\AW\D]G\>9P\^C\]V]GK\AlTVGZ@>9C\AGZ]CFGZ]CFG	Z]@GWl_\TZPlEVPG\AW\D]G\>9\FGCFG	\FG@GWl_\TZPlEVPG\AW\D]G\>9V]WP\^C\]V]G>9P\^C\]V]GWVP\WVAlKZ@>9C\AGZ]CFG	Z]@GWl_\TZPlEVPG\A W\D]G\>9\FGCFG	\FG@GWl_\TZPlEVPG\AW\D]G\>9V]WP\^C\]V]G>9QVTZ]>9	WVP\WVAlKC\AG^RCZ]CFGlWVP\WVA>9	WVP\WVAlKC\AG^RCZ]CFGlWVP\WVA>9	K\AlTVGC\AG^RCWVP\WVAK\AxVJ\FGCFG>9 	K\AlTVGC\AG^RCWVP\WVAK\AxVJ\FGCFG>9>9V]WqV[REZ\AR_