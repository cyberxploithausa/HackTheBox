NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNniNNC
C CCC
niNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNni
C
XniC
M<
 <RRUWMXnini
C<C
niCCCCK
RO
QCYC
C<
 < KRVCCSJXniCCCCCCCCCYCC<
 < KRVCCSJJXniCCCCC<Xnini 
 C!
CC<C
ni
niCCCCC_^C
RCC
QXniC!
XniniNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNniNNC C CC CWRUniNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNni
C
XniC
M<
 <RRUWMXnini
C <WRUC
niCCCCK
CYC
C<
 < KPCCSJXniCCCCCCCCCYCC<
 < KRVCCSJJXniCCCCC <WRUXnini 
 C!
CC <WRUC
ni
niCCCC K
JniCCCC
niCCCCCCCC C
C
niCCCCCCCCCCCCCASSSSAC^]CC_^CASSSSSSSSSSSSSSSRAXniCCCCCCCCCCCCCASSSRAC^]CC_^CASSSSSSSSSSSSSSRSAXniCCCCCCCCCCCCCASSRSAC^]CC_^CASSSSSSSSSSSSSRSSAXniCCCCCCCCCCCCCASSRRAC^]CC_^CASSSSSSSSSSSSRSSSAXniCCCCCCCCCCCCCASRSSAC^]CC_^CASSSSSSSSSSSRSSSSAXniCCCCCCCCCCCCCASRSRAC^]CC_^CASSSSSSSSSSRSSSSSAXniCCCCCCCCCCCCCASRRSAC^]CC_^CASSSSSSSSSRSSSSSSAXniCCCCCCCCCCCCCASRRRAC^]CC_^CASSSSSSSSRSSSSSSSAXniCCCCCCCCCCCCCARSSSAC^]CC_^CASSSSSSSRSSSSSSSSAXniCCCCCCCCCCCCCARSSRAC^]CC_^CASSSSSSRSSSSSSSSSAXniCCCCCCCCCCCCCARSRSAC^]CC_^CASSSSSRSSSSSSSSSSAXniCCCCCCCCCCCCCARSRRAC^]CC_^CASSSSRSSSSSSSSSSSAXniCCCCCCCCCCCCCARRSSAC^]CC_^CASSSRSSSSSSSSSSSSAXniCCCCCCCCCCCCCARRSRAC^]CC_^CASSRSSSSSSSSSSSSSAXniCCCCCCCCCCCCCARRRSAC^]CC_^CASRSSSSSSSSSSSSSSAXniCCCCCCCCCCCCCARRRRAC^]CC_^CARSSSSSSSSSSSSSSSAXniCCCCCCCCCCCCCC^]CC_^CASSSSSSSSSSSSSSSSAXniCCCCCCCCC XniCCCCC XniC!
XniniNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNniNNC
C niNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNni
C
XniC
M<
 <RRUWMXnini
C
C
niCCCCK
<RO
<QCYC
C<
 < KPCCSJXniCCCCCCCC(CYC
C<
 < KRVCCSJXniCCCCCCCCROQCYCC<
 < KRVCCSJJXniCCCCC
Xnini 
 C!
CC
C
niniCCCC
C RO QYC<
 < KRVCCSJXniCCCC C<C
niCCCCCCCCK
RO
QCYC
C<
 < KRVCCSJXniCCCCCCCCCCCCCYCC<
 < KRVCCSJJXniCCCCCCCCC XniCCCC C <WRUC
niCCCCCCCCK
CYC
C<
 < KPCCSJXniCCCCCCCCCCCCCYCC<
 < KRVCCSJJXniCCCCCCCCC XniCCCCCCCCCCCC
niCCCCCCCCCCCCCCCC/SCYC <WRUCCK
<RO RJXniCCCCCCCCCCCCCCCC/RCYC <WRUCCK
<QO QJXniCCCCCCCCCCCCCCCC/QCYC<CCK RO(ORJXniCCCCCCCCCCCCCCCC/PCYC<CCK QO(OQJXniniCCCCCCCCC!
X