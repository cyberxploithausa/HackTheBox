:::::::::::::::::9:7U~AdG7Px^g\yVyG7UxA7KxA7\gVeRcZx]9:::::::::::::::::9{ZuAvAn~VrV,>FdV7ZrVrdGsl{\pZtl&!9R{_,>>VyG~Gno\elpVc~@977g\eG?ZyCbG&~]gFc7	7ZydGsl{\pZtlaVtGxA?"s\`]c\7>97777xFcCbG7	7\bG7@cWH_xT~PHErPc\e&7WxDyGx'>977r]so\elpVc99vAt[~GrPcFeV7qr[vE~\eR{xU7KxAHTrG7Zd>QrT~]977xFcCbG7*~]gFc7KxA7ZyCbG%9r]sUVRaZxAv_,>>:::::::::::::::::>:dVt\yW7Px^g\yVyG7UxA7WrPxWrA7o!>:::::::::::::::::>_~QeReJ7ZrVr9b@r~VrV9@cWH_xT~PH&#v_{99r]cZcJ7WrPxWrAHo!~@977g\eG?ZyCbG7	7ZydGsl{\pZtlaVtGxA? 7WxDyGx',>7777\bGgFc-xFcdGsl{\pZtlaVtGxA?"s\`]c\7>,>77VyW7WrPxWrAHo!99vAt[~GrPcFeV7qr[vE~\eR{xU7WrPxWrAHo!~@9uVpZy>77Ce\tVd@?ZyCbG>>77QrT~]97777tRdV7ZyCbG7Zd>777777DVy5''7)xFcCbG7*5'''''''&,>777777DVy5'&7)xFcCbG7*5'''''''',>777777DVy5''7)xFcCbG7*5''''''&',>777777DVy5'&7)xFcCbG7*5'''''''',>777777DVy5&'7)xFcCbG7*5'''''&'',>777777DVy5&&7)xFcCbG7*5'''''''',>777777DVy5&'7)xFcCbG7*5''''&''',>777777DVy5&&7)xFcCbG7*5'''''''',>777777DVy5''7)xFcCbG7*5'''&'''',>777777DVy5'&7)xFcCbG7*5'''''''',>777777DVy5''7)xFcCbG7*5''&''''',>777777DVy5'&7)xFcCbG7*5'''''''',>777777DVy5&'7)xFcCbG7*5'&'''''',>777777DVy5&&7)xFcCbG7*5'''''''',>777777DVy5&'7)xFcCbG7*5&''''''',>777777DVy5&&7)xFcCbG7*5'''''''',>777777DVyxGVe@7)xFcCbG7*5'''''''',>7777VyW7Pv@r977r]sgAxPr@d9r]sUVRaZxAv_,>>:::::::::::::::::>:zR~]7Px^g\yVyG9:::::::::::::::::9{ZuAvAn~VrV,>FdV7ZrVrdGsl{\pZtl&!9R{_,>>VyG~GnzR~]7Zd>77CxAc~]gFcl&~]gFcl%-~]7@cWH_xT~PHErPc\e$s\`]c\7>97777o\exrJ7	7ZydGsl{\pZtlaVtGxA?"s\`]c\7>97777xFcCbG&xFcCbG%-xFcdGsl{\pZtlaVtGxA?"s\`]c\7>,>77VyW7^vZy99vAt[~GrPcFeV7qr[vE~\eR{xU7^vZy~@9977dZp]v_7WrPxWrA&sVt\sVe-dGsl{\pZtlaVtGxA?"s\`]c\7>977t\zCx]r]co\elpVc~@97777g\eG?ZyCbG&~]gFc7	7ZydGsl{\pZtlaVtGxA?"s\`]c\7>9777777xFcCbG7	7\bG7@cWH_xT~PHErPc\e&7WxDyGx'>97777r]st\zCx]r]c977t\zCx]r]csVt\sVel#K&7Zd>7777CxAc~]gFc-~]7@cWH_xT~PHErPc\e$s\`]c\7>9777777xFcCbG7	7\bG7@cWH_xT~PHErPc\e&7WxDyGx'>97777r]st\zCx]r]c9777777uVpZy>77777777'-sVt\sVel#K&7CxAczRg~]gFcl&sVt\sVe>977777777[7	7WrPxWrAHo!g\eG7^vC?ZyCbGH;WrPxWrA%,>77777777%-o\elpVcg\eG7^vC?WrPxWrA&o\exrJ;\bGgFc>977777777[ 7	7KxAHTrG7CxAczRgsVt\sVe;KxA\VnxFcCbG%,>>7777VyW7qr[vE~\eR{