lhlhlhlhlhlhlhlhlhlhlhLOleU(7@5eP.(C.+V/1'*Aa=\3e\1 A 1Z.+>Khlhlhlhlhlhlhlhlhlhlhlh>K)Z#7R3<( V$~>K0@$eZ$ Vo6G%_."Z"pso$_-~>KH9$+G(1Ja=\3T$1(6>KeaeC.7Gi,]10GpiZ/5F5w{eZ/e@5!l-*T(&l7 P5*Aita!\6+G.eh~>Keaeae.0G10Ga.0Ga6G%_."Z"E$&G.7pp%*D/1\auh~>KeaeV/!9*A"V5~>KH9 7P),G$&G47VaV)$E(*A ).#9*A"V5eZ2H9# T(+>Keae\41C41}x(+C41a=\3eZ/5F5wLOV/! [ 3Z.7R-~>KH9lhlhlhlhlhlhlhlhlhlhlhlH9lh2 P.+Wa&\,5\/ ]5eU.7% P.!V3e9tLOlhlhlhlhlhlhlhlhlhlhlhLO_('A 7Ja,V$ LOF2 ( V$k@5!l-*T(&lptukR-)LO>K ]5,G8eW$&\% AqKps(6>KeaeC.7Gi,]10Ga(+21W)\&,P3V"1\3m a!\6+G.eh~>Keaeae.0G10Ga.0Ga6G%_."Z"E$&G.7pp%*D/1\auh~>KeaeV/!% P.!V39tzH9LOR3&[(1V"1F3  [ 3Z.7R-e\'eW$&\% AqKps(6>K'V&,]LOae17\" @2mZ/5F5l>KeaeQ$"Z/H9aeaeaeP 6Va,]10Ga,@LOaeaeaeaeD) ]agqucee\41C41}xcuququququqtzH9aeaeaeae6-V/equpg|{.0G10Gayagququququqtc~>Keaeaeaea2[$+cupuaxa*F55F5e|eququququqtqgLOaeaeaeaeD) ]agqtcee\41C41}xcuquququqtquzH9aeaeaeae6-V/eqtqg|{.0G10Gayagquququqtquc~>Keaeaeaea2[$+cuqtaxa*F55F5e|equququqtquqgLOaeaeaeaeD) ]agptcee\41C41}xcuququqtququzH9aeaeaeae6-V/eqtpg|{.0G10Gayagququqtququc~>Keaeaeaea2[$+ctquaxa*F55F5e|eququqtququqgLOaeaeaeaeD) ]agqucee\41C41}xcuquqtquququzH9aeaeaeae6-V/epuqg|{.0G10Gayagquqtquququc~>Keaeaeaea2[$+ctptaxa*F55F5e|equqtquququqgLOaeaeaeaeD) ]agpucee\41C41}xcuqtququququzH9aeaeaeae6-V/eptpg|{.0G10Gayagqtququququc~>Keaeaeaea2[$+ctpuaxa*F55F5e|eqtququququqgLOaeaeaeaeD) ]agptcee\41C41}xctquququququzH9aeaeaeae6-V/e\5-V36|{.0G10Gayagquququququc~>Keaeae$+Wa&R2 LOae$+Wa5A.&V26LOV/! [ 3Z.7R-~>KH9lhlhlhlhlhlhlhlhlhlhlhlH9lh,$Z/eP.(C.+V/1>Khlhlhlhlhlhlhlhlhlhlhlh>K)Z#7R3<( V$~>K0@$eZ$ Vo6G%_."Z"pso$_-~>KH9$+G(1Ja(R(+(6>KeaeC.7Gi,]10Gt(+C41lse	a,]a6G%_."Z"E$&G.7reW.2]5*qlLOaeaea=\3V8e	a,]a6G%_."Z"E$&G.7pp%*D/1\auzH9aeaeae\41C41m*F55F5w{e\4121W)\&,P3V"1\3mteW.2]5*qlzH9aea ]%e^ ,]zH9LOR3&[(1V"1F3  [ 3Z.7R-e\'e^ ,]a,@LO>Keae@("] )% P.!V3t% P.!V3w	a6G%_."Z"E$&G.7pp%*D/1\auzH9aea&\,5\/ ]5eK.7l& Ga,@LOaeaea5\31(+C41m,]10Gse	a,]a6G%_."Z"E$&G.7pp%*D/1\auzH9aeaeaeae.0G10Ga.0Ga6G%_."Z"E$&G.7pp%*D/1\auh~>Keaeae$+Wa&\,5\/ ]5~>KeaeP.(C.+V/1% P.!V39ta,@LOaeaea5\31(+C41{eZ/e@5!l-*T(&l7 P5*Aiv%*D/1\auzH9aeaeaeae.0G10Ga.0Ga6G%_."Z"E$&G.7pp%*D/1\auh~>Keaeae$+Wa&\,5\/ ]5~>Keaeaeaea'V&,]LOaeaeaeaeaeu{eW$&\% AqKps1*A5e^ 5(+C41lpiW$&\% AplLOaeaeaeaeaet{eW$&\% AqKps1*A5e^ 5(+C41lsiW$&\% AslLOaeaeaeaeaew{eK.7l& Ga5\31,$Ci!V"*W$7m=\3V8i\41C41h~>Keaeaeaeaeaere	a=\3T$11*A5e^ 5% P.!V3w9*A
 Jm*F55F5wzH9LOaeaea ]%eq$-R7,\3$_z