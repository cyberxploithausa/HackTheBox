NyNyNyNyNyNyNyNyNyNyNyNyNyNyNyNyNyn^NyC2
& C79;1 C2&C,&C;15=:n^NyNyNyNyNyNyNyNyNyNyNyNyNyNyNyNyNyn^=&&t
11XYi!1C=1z ;= ReU`M58XYiYi1 
 t;1t
'n^CtCt; K=$ Rx
:!fCnC=t ;= 1  &KeVt;:;CdJon^CtCtCtCt!$ CnC; C'0<83
7<"7;|RaC0# tS}Jon^CtCt:t;1on^n^& <
 7!1C<"
;5t2C,&<3 C=Yi63
:n^CtCt!$ Ch^t
:!eC,&C=$ Qon^:t!15=&8XYiYiyNyNyNyNyNyNyNyNyNyNyNyNyNyNyNyNyNYiyNt1 ;0C79;1 C2&C070&C`eUYiyNyNyNyNyNyNyNyNyNyNyNyNyNyNyNyNyNYi8
65-C=1on^'t
11M'0<83
7<eRbWz8on^n^:=-C070&<`eUt
'n^CtCt; K=$ CnC=t ;= 1  &KgC0# tS}XYitCtCtCtC; !tYt!t ;= 1  &KeVt;:;CdJ}XYitCtC10C070&<`eUon^n^& <
 7!1C<"
;5t2C070&<`eUt
'n^1=YitCtC$; 1'K=$ JYitCtC63
:n^CtCtCtCt 51C=$ C=YitCtCtCtCtCtC#1tAdSdSvCi]t!$ Ch^tAdSdSdSdSdSdSdSdRvXYitCtCtCtCtCtC#1tAdSdRvCi]t!$ Ch^tAdSdSdSdSdSdSdSeSvXYitCtCtCtCtCtC#1tAdSeSvCi]t!$ Ch^tAdSdSdSdSdSdSdRdSvXYitCtCtCtCtCtC#1tAdSeRvCi]t!$ Ch^tAdSdSdSdSdSdSeSdSvXYitCtCtCtCtCtC#1tAdRdSvCi]t!$ Ch^tAdSdSdSdSdSdRdSdSvXYitCtCtCtCtCtC#1tAdRdRvCi]t!$ Ch^tAdSdSdSdSdSeSdSdSvXYitCtCtCtCtCtC#1tAdReSvCi]t!$ Ch^tAdSdSdSdSdRdSdSdSvXYitCtCtCtCtCtC#1tAdReRvCi]t!$ Ch^tAdSdSdSdSeSdSdSdSvXYitCtCtCtCtCtC#1tAeSdSvCi]t!$ Ch^tAdSdSdSdRdSdSdSdSvXYitCtCtCtCtCtC#1tAeSdRvCi]t!$ Ch^tAdSdSdSeSdSdSdSdSvXYitCtCtCtCtCtC#1tAeSeSvCi]t!$ Ch^tAdSdSdRdSdSdSdSdSvXYitCtCtCtCtCtC#1tAeSeRvCi]t!$ Ch^tAdSdSeSdSdSdSdSdSvXYitCtCtCtCtCtC#1tAeRdSvCi]t!$ Ch^tAdSdRdSdSdSdSdSdSvXYitCtCtCtCtCtC#1tAeRdRvCi]t!$ Ch^tAdSeSdSdSdSdSdSdSvXYitCtCtCtCtCtC#1tAeReSvCi]t!$ Ch^tAdRdSdSdSdSdSdSdSvXYitCtCtCtCtCtC#1tAeReRvCi]t!$ Ch^tAeSdSdSdSdSdSdSdSvXYitCtCtCtCtCtC#1t 1'Ci]t!$ Ch^tAdSdSdSdSdSdSdSdSvXYitCtCtCtC10C7'on^CtCt:t&7'on^:t!15=&8XYiYiyNyNyNyNyNyNyNyNyNyNyNyNyNyNyNyNyNYiyNt5
:C79;1 n^NyNyNyNyNyNyNyNyNyNyNyNyNyNyNyNyNyn^=&&t
11XYi!1C=1z ;= ReU`M58XYiYi1 
 t5
:C=YitCtC$&|
:!Rx
:!QtYt
:C'0<83
7<"7;|Pt;:;CdJon^CtCtCtCt;-CnC=t ;= 1  &KeVt;:;CdJon^CtCtCtCt!$ Rx!$ QtYt!t ;= 1  &KeVt;:;CdJ}XYitCtC10C9=on^n^& <
 7!1C<"
;5t2C9=t
'n^n^CtCt=:8C070&Rx1 ;1fYt ;= 1  &KeVt;:;CdJon^CtCt ;$::t;1t
'n^CtCtCtCt; K=$ Rx
:!fCnC=t ;= 1  &KeVt;:;CdJon^CtCtCtCtCtCt!$ CnC; C'0<83
7<"7;|RaC0# tS}Jon^CtCtCtCt:t ;$::on^CtCt ;$::t1 ;1W,RbC=YitCtCtCtC$&|
:!tYt
:C'0<83
7<"7;|Pt;:;CdJon^CtCtCtCtCtCt!$ CnC; C'0<83
7<"7;|RaC0# tS}Jon^CtCtCtCt:t ;$::on^CtCtCtCtCtCt1=YitCtCtCtCtCtCtCtCStYt1 ;1W,RbC$&t5|
:!Rx1 ;1eJon^CtCtCtCtCtCtCtCt/eCnC070&<`eUt; C9$K=$ <fO070&Q}XYitCtCtCtCtCtCtCtCQtYt;1t; C9$K070&Rx;-O; !eJon^CtCtCtCtCtCtCtCt/gCnC,&<3 C$&t5|1 ;1fO,&(1x!$ Q}XYiYitCtCtCtC10C<"
;5o